--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   00:34:20 05/19/2023
-- Design Name:   
-- Module Name:   /home/ise/Documents/ContadorHorasProj/tb_contadorHoras.vhd
-- Project Name:  ContadorHorasProj
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: ContadorHoras
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_contadorHoras IS
END tb_contadorHoras;
 
ARCHITECTURE behavior OF tb_contadorHoras IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT ContadorHoras
    PORT(
         CLK : IN  std_logic;
         RST : IN  std_logic;
			LAP_ENABLE : IN  std_logic;
         LAP : OUT  std_logic;
         OUTPUT : OUT  std_logic_vector(7 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal CLK : std_logic := '0';
   signal RST : std_logic := '0';
   signal LAP_ENABLE : std_logic := '1';
	
 	--Outputs
   signal LAP : std_logic;
   signal OUTPUT : std_logic_vector(7 downto 0);

   -- Clock period definitions
   constant CLK_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: ContadorHoras PORT MAP (
          CLK => CLK,
          RST => RST,
          LAP => LAP,
			 LAP_ENABLE => LAP_ENABLE,
          OUTPUT => OUTPUT
        );

   -- Clock process definitions
   CLK_process :process
   begin
		CLK <= '0';
		wait for CLK_period/2;
		CLK <= '1';
		wait for CLK_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      wait;
   end process;

END;
